`define FTIME 30000000
module tb_testbench();
reg CLK, RESETB;
reg [7:0] DATA;
wire [12543:0] OUTPUT;
wire VALID;
integer fp;

cnn c1(
    .axi_clk(CLK),
    .axi_rst_n(RESETB),
    .i_data_valid(1'b1),
    .i_data(DATA),
    .o_data_valid(VALID),
    .o_convoledData(OUTPUT) //32*7*7*8
);


initial begin
    CLK     = 1'b0;
    RESETB  = 1'b0;
    #10 fp = $fopen("output.txt", "w");
    #`FTIME;
    $fclose(fp);
    $finish;
end


// test condition
initial begin
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00011111 ;
#100 DATA = 00101000 ;
#100 DATA = 10000001 ;
#100 DATA = 11101010 ;
#100 DATA = 11101010 ;
#100 DATA = 10011111 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 01000100 ;
#100 DATA = 10010110 ;
#100 DATA = 11101111 ;
#100 DATA = 11111110 ;
#100 DATA = 11111101 ;
#100 DATA = 11111101 ;
#100 DATA = 11111101 ;
#100 DATA = 11010111 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 10011100 ;
#100 DATA = 11001001 ;
#100 DATA = 11111110 ;
#100 DATA = 11111110 ;
#100 DATA = 11111110 ;
#100 DATA = 11110001 ;
#100 DATA = 10010110 ;
#100 DATA = 01100010 ;
#100 DATA = 00001000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00010011 ;
#100 DATA = 10011010 ;
#100 DATA = 11111110 ;
#100 DATA = 11101100 ;
#100 DATA = 11001011 ;
#100 DATA = 01010011 ;
#100 DATA = 00100111 ;
#100 DATA = 00011110 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 10010000 ;
#100 DATA = 11111101 ;
#100 DATA = 10010001 ;
#100 DATA = 00001100 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00001010 ;
#100 DATA = 10000001 ;
#100 DATA = 11011110 ;
#100 DATA = 01001110 ;
#100 DATA = 01001111 ;
#100 DATA = 00001000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 10000110 ;
#100 DATA = 11111101 ;
#100 DATA = 10100111 ;
#100 DATA = 00001000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 11111111 ;
#100 DATA = 11111110 ;
#100 DATA = 01001110 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 11001001 ;
#100 DATA = 11111101 ;
#100 DATA = 11100010 ;
#100 DATA = 01000101 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00110111 ;
#100 DATA = 00000110 ;
#100 DATA = 00000000 ;
#100 DATA = 00010010 ;
#100 DATA = 10000000 ;
#100 DATA = 11111101 ;
#100 DATA = 11110001 ;
#100 DATA = 00101001 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00011001 ;
#100 DATA = 11001101 ;
#100 DATA = 11101011 ;
#100 DATA = 01011100 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00010100 ;
#100 DATA = 11111101 ;
#100 DATA = 11111101 ;
#100 DATA = 00111010 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 11100111 ;
#100 DATA = 11110101 ;
#100 DATA = 01101100 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 10000100 ;
#100 DATA = 11111101 ;
#100 DATA = 10111001 ;
#100 DATA = 00001110 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 01111001 ;
#100 DATA = 11110101 ;
#100 DATA = 11111110 ;
#100 DATA = 11111110 ;
#100 DATA = 11111110 ;
#100 DATA = 11011001 ;
#100 DATA = 11111110 ;
#100 DATA = 11011111 ;
#100 DATA = 00110010 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 01110100 ;
#100 DATA = 10100101 ;
#100 DATA = 11101001 ;
#100 DATA = 11101001 ;
#100 DATA = 11101010 ;
#100 DATA = 10110100 ;
#100 DATA = 00100111 ;
#100 DATA = 00000011 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#100 DATA = 00000000 ;
#10 $fwrite(fp, "%b\n",OUTPUT);
end

always begin
    #50 CLK = ~CLK; // 100ns period pulse
end

initial begin
    $dumpfile("tb_testbench_out.vcd");
    $dumpvars(0, tb_testbench);  
end

endmodule


// ref by https://github.com/vipinkmenon
module cnn #(
    parameter F = 28, // feature
    parameter B = 8 // bit size
)(
    input axi_clk,
    input axi_rst_n,
    // slave i/f
    input i_data_valid,
    input [B-1:0] i_data,
    // output o_data_ready,
    // master i/f
    output [15:0] o_data_valid,
    // output [B-1:0] o_data,
    // input i_data_ready,
    // interrupt
    output o_intr,
    output [16*B-1:0] o_convoledData //32*7*7*8
);

    wire [3*3*B-1:0] pixel_data_conv1;
    wire pixel_data_conv1_valid;

    wire [16*3*3*B-1:0] pixel_data_conv2;
    wire [15:0] pixel_data_conv2_valid;

    wire [255:0] convoled_data_conv2;
    wire [31:0] convoled_data_conv2_valid;

    wire axis_prog_full;
    wire [16*B-1:0] L1_convoled_data;
    wire [16-1:0] L1_convoled_data_valid;

    reg [16*B-1:0] conv1_bias;
    reg [1151:0] conv1_weight;
    //reg [255:0] conv2_bias;
    //reg [36863:0] conv2_weight;

    wire intr_L1;
    assign o_intr = intr_L1;
    //wire [15:0] intr_L2;
    
    // assign o_data_ready = !axis_prog_full;// if buffer full, it means not ready to get data

    // assign valid = i_data_valid[0]
    
    wire [B-1:0] data;
    assign data = intrCnt<=F-3 ? i_data : 'b0;
    wire inputValid;
    wire paddingValid;
    assign inputValid = i_data_valid | paddingValid; // >> 벨리드 28클럭 유지해서 0 두줄 넣도록 하는 부분 추가구현 필요

    reg [$clog2(F)-1:0] intrCnt;
    always@(posedge axi_clk)begin
        if(!axi_rst_n | (intrCnt==(F-1)) | (intrCnt==(F-2) & lineCnt==F))
            intrCnt <= 0;
        else if(intr_L1)
            intrCnt <= intrCnt + 1;
    end

    assign paddingValid = intrCnt>F-4 & lineCnt != F;
    
    reg [$clog2(F+1)-1:0] lineCnt;
    always@(posedge axi_clk)begin
        if(!axi_rst_n | lineCnt == F)
            lineCnt <= 0;
        else if(intrCnt == F-3 | intrCnt == F-2)begin
            lineCnt <= lineCnt + 1;
        end
    end

    ctrl L1_ctrl(
        .i_clk(axi_clk),
        .i_rst(!axi_rst_n),
        .i_pixel_data(data),
        .i_pixel_data_valid(inputValid),
        .o_pixel_data(pixel_data_conv1),
        .o_pixel_data_valid(pixel_data_conv1_valid),
        .o_intr(intr_L1)
    );

    conv_L1 L1(
        .i_clk(axi_clk),
        .i_pixel_data(pixel_data_conv1),
        .i_pixel_data_valid(pixel_data_conv1_valid),
        .i_weight(conv1_weight),
        .i_bias(conv1_bias),
        .o_convloed_data(L1_convoled_data),
        .o_convloed_valid(L1_convoled_data_valid)
    );


    // ctrlL2 L2_ctrl(
    //     .i_clk(axi_clk),
    //     .i_rst(!axi_rst_n),
    //     .i_pixel_data(L1_convoled_data),
    //     .i_pixel_data_valid(L1_convoled_data_valid),
    //     .i_weight(conv2_weight),
    //     .i_bias(conv2_bias),
    //     .o_pixel_data(pixel_data_conv2),
    //     .o_pixel_data_valid(pixel_data_conv2_valid),
    //     .o_intr(intr_L2)
    // );

    // conv_L2 L2(
    //     .i_clk(axi_clk),
    //     .i_convloed_data(pixel_data_conv2[j]),
    //     .i_convloed_valid(pixel_data_conv2_valid[j]),
    //     .o_convloed_data(convoled_data_conv2),//[32*8-1:0] == [255:0]
    //     .o_convloed_valid(convoled_data_conv2_valid)
    // );



    // reg [$clog2(49)-1:0] outIdx;
    // always@(posedge axi_clk)begin
    //     if(axi_rst_n)
    //         outIdx <= 'd0;
    //     else if(convoled_data_conv2_valid)begin
    //         if(outIdx <'d48)
    //             outIdx <= outIdx+1;
    //         else
    //             outIdx <= 0;
    //     end
    // end

    // reg [12543:0] outBuff;
    // always@(posedge axi_clk)begin
    //     if(axi_rst_n)
    //         outIdx <= 'd0;
    //     else
    //         outBuff[outIdx*256+:256] <= convoled_data_conv2;
    // end

    assign o_convoledData = L1_convoled_data;
    assign o_data_valid = L1_convoled_data_valid;
    // assign o_intr = intr_L1 ||  (|intr_L2);

    initial begin
        conv1_bias[7:0] <= 8'b01111011; //normalized bias=123.0000
        conv1_weight[71:0] <= 72'b10100000_10010011_10000001_10011011_10011001_01100011_01100111_10001100_10000001;
        conv1_bias[15:8] <= 8'b01111010; //normalized bias=122.0000
        conv1_weight[143:72] <= 72'b10100000_10010101_10000101_01110111_10010100_01011100_10010001_10000011_01111111;
        conv1_bias[23:16] <= 8'b01111111; //normalized bias=127.0000
        conv1_weight[215:144] <= 72'b10100000_10001110_10001100_10001110_10101000_10100001_10010110_10001110_10000100;
        conv1_bias[31:24] <= 8'b01111101; //normalized bias=125.0000
        conv1_weight[287:216] <= 72'b01100101_01011001_01111010_10001001_10101101_01111111_10000100_01101111_01011110;
        conv1_bias[39:32] <= 8'b01101110; //normalized bias=110.0000
        conv1_weight[359:288] <= 72'b01110010_10101110_01100101_01100010_10001110_10001100_01101000_10000010_10001110;
        conv1_bias[47:40] <= 8'b01110111; //normalized bias=119.0000
        conv1_weight[431:360] <= 72'b01110011_10001111_10011100_10001000_10111100_10110000_01111000_01110101_01110100;
        conv1_bias[55:48] <= 8'b01111011; //normalized bias=123.0000
        conv1_weight[503:432] <= 72'b01100001_10000011_01110111_10100001_01111010_01111000_10000110_01100101_01110110;
        conv1_bias[63:56] <= 8'b01111101; //normalized bias=125.0000
        conv1_weight[575:504] <= 72'b01110001_10000010_10011111_01110011_01101011_10001011_01101000_01101010_01111010;
        conv1_bias[71:64] <= 8'b01111111; //normalized bias=127.0000
        conv1_weight[647:576] <= 72'b10001111_10100100_10010011_10011111_10010000_10010000_01110010_01110100_01101011;
        conv1_bias[79:72] <= 8'b01111110; //normalized bias=126.0000
        conv1_weight[719:648] <= 72'b01010100_10100100_10100001_01110000_01110101_01110101_01100000_01111100_10000100;
        conv1_bias[87:80] <= 8'b01111010; //normalized bias=122.0000
        conv1_weight[791:720] <= 72'b01101000_01100001_10010010_01111100_01111111_10010110_01111100_01101010_01101000;
        conv1_bias[95:88] <= 8'b01101110; //normalized bias=110.0000
        conv1_weight[863:792] <= 72'b10010010_01110101_10000010_01101110_01111011_01101000_01111001_10001011_01111010;
        conv1_bias[103:96] <= 8'b01110111; //normalized bias=119.0000
        conv1_weight[935:864] <= 72'b01111111_01110110_10000001_01110001_01101111_01111011_10000001_10000101_01111100;
        conv1_bias[111:104] <= 8'b01110111; //normalized bias=119.0000
        conv1_weight[1007:936] <= 72'b10000000_01111011_01011100_01111100_01010110_01111011_10100000_10000010_10000010;
        conv1_bias[119:112] <= 8'b01111101; //normalized bias=125.0000
        conv1_weight[1079:1008] <= 72'b10010100_10011111_10010110_10100010_10101111_10100001_10010000_10001000_10001101;
        conv1_bias[127:120] <= 8'b01111010; //normalized bias=122.0000
        conv1_weight[1151:1080] <= 72'b01111101_01111011_01111110_01111001_01110111_01110010_10000100_01110110_01111000;
    end
    
    // initial begin
    //     conv2_bias[7:0] <= 8'b01100000; //normalized bias=96.0000
    //     conv2_weight[1151:0] <= 1152'b01101101_10101101_10001110_10101001_11000101_01111010_01100001_01101100_01110001_01111010_01111011_01111101_01101101_10000110_10001001_10010010_01111000_10001000_10001011_10000001_01101101_01110000_01110010_01111000_01110111_01111101_10000000_01111101_01111101_01111101_10010100_10000101_01110111_01100001_10001010_01111001_01111011_10010010_01111100_01111011_01110011_10000000_01111111_01111011_10001001_01111100_10000001_10010110_01100100_01110100_01111100_01110111_01110111_10000001_01111111_10010100_01111110_01110010_10000010_10001110_01111101_01111001_01101111_01111010_10001001_01110011_01101110_01110010_01110011_10011010_01100101_01111111_10000101_10001011_01110111_10010010_10010110_10000100_10000000_01101111_10001000_01110010_01101110_10000110_10000010_10000110_10010100_01111111_01111101_01110110_01110110_01111101_10000110_01110000_10010010_01110011_01101111_01111101_01110011_01111111_01110101_10001111_10001000_10010011_01110110_01111100_10000101_01101001_10000000_01110100_01110000_10001110_01111011_01111111_10000001_01111110_01111000_10010000_01111100_01100110_01111110_10000110_10000100_01111101_10000110_10010010_10010001_01101001_01111000_10000100_10010001_10000001_01110111_01111111_01111110_01111001_10001101_01111011_01110111_10010000_01111001_10000010_01111100_01111100;
    //     conv2_bias[15:8] <= 8'b10000001; //normalized bias=129.0000
    //     conv2_weight[2303:1152] <= 1152'b10001010_10010110_10101000_01001010_00111111_01011110_10100111_10000110_01111111_10000111_01110010_01111011_10010101_10010001_10000100_10000001_01111101_10001101_01111100_01111101_01110110_10001011_01100000_10000100_10011001_01101101_10000111_10000101_10011001_01101101_01100001_10001000_01110110_10000001_01111010_01100110_01111111_01111001_10000101_01110010_10001101_10000000_10000011_01110111_01100110_10000010_10000001_10001001_10000010_01111011_01100101_01110011_01111111_01110111_10000000_01101011_10010010_10001001_10000010_01111100_01111010_01110111_01110000_01111110_10000100_10000111_01111100_01110110_10010010_10000101_10000101_01101110_10001111_10001101_01100110_10010001_10001010_01100000_01101000_10000010_01110101_01111110_01110000_10010001_01110111_10001101_01100111_10000010_10000100_10001000_10001011_10000100_01111011_10000011_10000100_10000010_10010100_01110110_01111000_01110110_10010010_01111111_01110101_10001001_01110111_01111111_10001110_01111110_01011011_01110001_10000111_01111100_10000001_10010001_01111101_01111100_10000001_01011110_10000111_10001001_10010101_01110101_01111011_10001111_10000111_10001101_10001001_10001000_01110100_10001001_01111011_01111000_10000101_10000011_10000000_10000010_10010111_01100100_01111101_01110100_10000010_10000001_01100010_10001100;
    //     conv2_bias[23:16] <= 8'b01011011; //normalized bias=91.0000
    //     conv2_weight[3455:2304] <= 1152'b10010110_00111010_00100000_10101011_11010011_10100000_01110001_10011001_10010100_10010101_10000010_10000001_01101111_01110100_01101110_10001011_10000011_01101101_01111011_01110010_01111101_01111111_10001110_01111101_10001111_01110000_01111100_01111001_01101101_10000000_10000111_10001100_01111111_10010000_01111001_10000101_01111011_01100100_10000010_10000000_10000111_10001110_10000111_01110100_10000010_01101000_01101110_01101101_10010110_10001101_01111111_01111111_01110110_01111010_10001001_10000011_01110001_01101101_10000010_01110010_10001010_10000110_10001010_10000001_10001000_01111101_01101011_01111101_01100011_10000001_10000101_01111101_01111100_01111010_01101010_10001010_01111000_01111001_10001010_10001101_01110110_10000100_10000100_01101101_10000111_01110100_01110101_01111001_10001110_10000011_10000110_10010000_10001001_01101010_10010000_01110100_01110100_01110001_01100000_10001001_10001011_01111101_10000101_10001001_01110100_10000111_10000000_10000010_01110001_01101101_01110011_10000000_01101111_10000101_01110011_10001100_10001100_10000000_10000011_10001100_01111011_10000000_01111101_10001001_10010010_01111010_01110011_10000011_10011000_01110100_01111000_01111111_10000000_10000000_10010111_01111101_01101001_01111010_10001011_10011011_01111101_10001010_01111011_10001100;
    //     conv2_bias[31:24] <= 8'b01110110; //normalized bias=118.0000
    //     conv2_weight[4607:3456] <= 1152'b10000110_01100101_01110110_01111010_10110011_10001010_01111101_10011001_01101001_10000000_01101011_01101111_10000110_10001010_10010001_01111110_01100001_01111010_01111111_01110100_01111010_10001001_01111111_01111010_01110100_10010100_01110111_10001000_01111100_01110001_10000010_10000001_10010000_10000110_10001011_10000110_10001100_01110110_01111011_01110101_10001010_10001001_10001011_10010011_01111001_01111000_01110011_01111010_10000100_01111111_01111011_01111000_10010101_10001100_10001010_10001000_01110111_10001100_01110101_10000001_10000010_10000001_01110101_10000001_01101011_01111011_10000101_10001010_10001011_10000101_01100110_10001010_01101110_10001111_01110010_10000100_10011001_01111101_01111010_01101111_10001010_01110001_10010100_01110101_01101010_10000001_01110001_01111100_10010101_01110101_10001011_01101001_10000001_10001000_10000100_10000001_10000010_01101000_10001000_01110011_01110011_01101110_10010011_01110111_01111111_01110000_01110001_10001000_01101011_01111011_10001010_10000010_01110111_01111101_01110001_10001000_10001010_01111010_01111000_10010010_01100011_10000111_01111011_10001001_10001001_01111101_01110001_01101111_01101111_10000011_01110110_01111111_01110001_01111011_10000000_01011111_10000100_10001011_01111000_01110101_01110101_01111101_10000010_01111110;
    //     conv2_bias[39:32] <= 8'b01111110; //normalized bias=126.0000
    //     conv2_weight[5759:4608] <= 1152'b01111100_10011100_01110111_01100011_01101110_01011011_01111011_10000000_01111101_01111010_10000101_01110110_01111110_01111010_10000011_10010100_10001011_01110111_10000010_10000000_01111001_10001100_01101010_10010000_01111010_10000110_10001101_10000100_10010010_10000101_01100011_01111100_10011000_01100010_10001100_01110010_10000101_10000000_01111101_01111000_01110100_10010000_10000011_01111111_01101110_10001110_01111100_01110011_10010111_01111010_10000000_01110001_10000010_01111101_01110000_10001001_10000110_01110100_10000001_10000000_10000100_10010001_01101110_10010010_10001011_10001000_01111100_01101110_10010000_10001101_10100100_10011100_01110111_10000101_01111000_10001000_10000110_01110001_10000000_10000110_10000110_01110111_10000001_01111111_10001001_01111011_10001010_10010001_01100010_01110000_10000111_01110100_01101000_01101010_10000010_10001000_01111100_01110010_01111111_10000001_10001111_01111011_01110000_10010001_01111100_01101111_01111111_01111110_01110001_01110001_01110100_10000000_01110001_10000101_01110001_01111100_10000110_01101110_01100011_01111100_01111011_10000000_10001011_10000001_01101100_01111011_10000010_10000011_01111100_10010101_10000010_01111001_01111001_10000100_01110100_10000110_01111011_10000100_10011111_01111011_01111111_01110101_10001000_01110110;
    //     conv2_bias[47:40] <= 8'b01111000; //normalized bias=120.0000
    //     conv2_weight[6911:5760] <= 1152'b10011010_01110011_01010000_10101110_01101111_01111000_10001001_01010011_01111001_10010101_10001001_10100001_10001000_10001110_01111101_01111110_01100011_10011011_10010100_10010110_01111010_01110001_01101010_01110110_01111110_01100001_10000100_10000010_01110010_10000100_10011010_01111101_01111001_10001110_01111010_01110110_01111011_01101010_01111101_01101100_10000111_01111010_10011010_01101100_10001011_10001000_10000000_10000010_10001100_10000110_01111000_10001110_01111010_01101111_01110110_10001100_10001101_10000011_01111011_01101010_10000111_10000011_01110000_01111101_10011100_10000001_01100101_10001011_01111001_01110000_01100111_01111010_01110000_10001111_01101010_10010101_10010001_01110011_10001011_01111110_01101110_01101011_01111100_01101011_01101101_01110111_10000010_10001011_10000000_01101101_10000100_10000011_01111010_10000010_10000000_10000000_01111110_10001000_10001010_01110110_10001001_10010011_10001010_10010111_10000001_10000111_01110010_10011011_01110110_10001010_10001010_10010110_01101100_10000011_01111101_01110101_01101100_01110011_10000011_01110100_10000001_01111101_01110011_01110101_10000010_01111011_10000100_10001000_01111001_01111111_01101110_10000100_10000100_10001111_10001101_10010101_01110100_01101000_10000001_01111101_10000010_10000010_10001101_10001110;
    //     conv2_bias[55:48] <= 8'b01111111; //normalized bias=127.0000
    //     conv2_weight[8063:6912] <= 1152'b10011110_10011110_10011000_01111110_10011010_01100111_00110001_00110010_00111011_10010001_10000111_10000000_10000001_01100101_10000101_01111110_01110010_01110100_10000100_01110100_01100010_01110101_01111111_01111100_10001111_01110010_10000101_01101110_01110010_01111110_01111101_01111100_10000111_10010111_10000011_10001101_01101110_10010011_10010000_01111000_10000100_10010011_01110001_10001000_01011100_10010010_01111101_10001000_10001101_01110100_01110101_01101000_01111101_01101111_01110110_01110000_10001111_10000111_01110010_10010001_10010001_10000100_10001101_01110010_01101011_01111001_01110010_10001110_01110110_10000111_10010100_01111011_10001000_10001000_01111110_01111111_10001001_01111001_10000101_01111000_01110100_01111111_01110000_10010001_01110101_10000010_01111000_10001100_01111001_10000010_10001010_01111110_01111110_01110101_01111000_10001001_01110101_10010111_01111011_01110111_10000011_01111000_01101110_10001000_01110011_01110011_01111001_01110111_01101111_01111010_01111110_01111111_10000111_01111001_10000110_10011100_01101111_01111011_01111010_10011000_10000111_01110100_10001000_10010100_01111110_01110101_10010001_10000001_01110111_01101110_01101111_10000111_10001000_01111100_10000101_10010000_10000001_10000110_10000100_10010100_01111110_01111000_10000000_10001001;
    //     conv2_bias[63:56] <= 8'b01001110; //normalized bias=78.0000
    //     conv2_weight[9215:8064] <= 1152'b01001010_10111110_01110000_00110001_11011000_01101111_01101000_10101011_01100110_10001010_10001111_01111000_01111010_10000111_10000010_10000011_10001000_01111011_01111110_01101101_01111100_10010000_10000111_10010100_01110000_01100000_01111111_10001101_10000001_01111011_10001100_10000010_10010010_01101011_01111001_01110101_10001101_10010100_10000101_01100101_10000101_01100101_10000110_01101100_10001001_10000100_01101101_01101101_01101111_01101011_01111111_01110000_01111001_01111110_01101111_10000011_01111001_10000001_10001101_01101111_10000100_01111111_10010001_01110000_10001010_01101010_01100000_01101000_10000101_01110001_10000001_10000000_10001010_10000111_01110110_01110000_01110111_10001101_10010000_01111100_01111010_10000100_10000010_10001100_10010110_01101111_01110110_01111110_01110111_01111110_10001111_10000010_10000111_10000000_01100011_10001101_01111000_01101011_01101000_01111000_10001010_01110011_10010001_10000010_10001000_01111001_10000110_10000101_10000011_01101011_01111000_01111100_01111111_10000011_01111000_10000011_10000110_10001001_10001001_01111101_01111000_01110110_10011001_01110010_01111101_10001100_10000110_10000010_10001010_01111011_10010001_10001000_01111101_10010000_01111010_10000000_10000100_01110010_10000111_10001100_10001110_10000001_01110111_10000111;
    //     conv2_bias[71:64] <= 8'b01111100; //normalized bias=124.0000
    //     conv2_weight[10367:9216] <= 1152'b01111010_10000100_01110101_01110100_01100001_10000100_01110000_10000001_01110101_10001011_01110101_01111101_10001110_10010010_10000100_01110010_10000000_01111100_01110001_10000000_01110111_10000100_10000101_10010000_10000100_01101110_10011001_10000110_01110011_01110011_10010000_01111011_10001001_01110010_10001111_10010000_10000010_10001101_10000010_10001010_10011000_10010001_01111100_01111101_10000010_10010001_01111001_01011111_10000011_01110110_01110101_10010011_01111001_10000001_01101100_10001001_01100111_10000001_10100000_01111110_01111000_10000011_10000011_01111001_10010101_01101110_10000010_10001000_01111011_01100010_10000000_01100010_01111000_01100011_10000111_01110010_10001111_10011000_01111100_10001011_10010100_10001011_01110110_10000110_10000011_01111101_01110101_01100110_10100011_10011011_10001110_10000011_10001000_10000101_01111010_10000000_01111010_10000010_01110111_01111100_01110010_10000100_10000010_01111001_10000000_01110111_10011100_01111001_01101111_10001111_01111011_01101011_01110111_10000001_01101011_01100110_01101001_10000011_10000010_10001011_01101101_10010100_10001001_10000011_01110110_10010111_01101011_01111110_01110011_10011000_10011011_10000001_10000101_01111101_10001101_01111010_10001110_01101111_10011011_01110100_10000010_01111011_01110111_01101100;
    //     conv2_bias[79:72] <= 8'b01110001; //normalized bias=113.0000
    //     conv2_weight[11519:10368] <= 1152'b10011111_01001010_01101100_11001000_01001100_01100110_10010010_00110110_10010000_01111111_01111001_10001011_10010010_01111001_01100101_10000100_10001001_01100111_10000010_01111100_01111110_01111110_10000001_10000110_10001001_10010000_10001010_10000000_10000010_01111011_10001101_01110100_10000011_01111110_01110000_10001101_01111111_10010010_01111101_01111001_10000100_10000000_10000011_01110101_01110000_01110000_10010010_10000110_10001111_01101011_10010110_10000001_01101110_01110010_01011010_10001000_01111010_01110100_10000000_01111111_10001110_01101110_01100111_10001111_01110000_10001101_01111100_01111001_10000111_01110001_10000011_01110101_01110111_01110011_01100000_10000000_01101001_10000001_01110000_10000111_01110100_10001011_01111110_01110100_10000101_10001010_01111000_01110100_01111100_10001011_10001011_01101010_10000110_01111101_01101110_10001101_10000000_01111100_10001000_10001001_01110011_01111110_01110011_10000101_01110000_01111110_01110011_01101011_10000101_10001010_01110010_01111110_10000001_01111001_10000010_10000001_10000001_01110011_10000111_10011000_10000111_01101101_10000011_10000010_01101010_01110001_01111100_10001000_01111010_01110001_01110101_10000101_01111100_01111111_10000010_10001111_01110111_10000111_01110111_01111101_10000011_10000110_10000001_10000000;
    //     conv2_bias[87:80] <= 8'b01111011; //normalized bias=123.0000
    //     conv2_weight[12671:11520] <= 1152'b01110100_01110011_01110111_01111010_01110001_01110011_10000000_01110001_01101111_10010001_01111100_01101011_01111100_01111011_10000111_01111000_01110011_10000001_01101111_10000100_01111000_10000011_10000110_01110010_01110110_10010101_01110110_10000100_01110010_10001010_01110001_01110101_10000100_01110100_01110110_10001100_10000010_01111111_10000011_01111101_10000111_10000011_01101010_01111000_01110011_01111101_10000000_10001100_10001001_10001000_01110100_10000101_01111100_10000011_01111101_10001000_01111011_01111101_01111010_01110010_01111101_01111111_01100000_01111100_10000000_10000010_10000100_10001011_01111010_01111001_01110100_01111101_10001001_10001000_01101111_10000101_01101001_01100100_10001001_10001010_10001010_10001010_01110101_01111101_01111010_10000001_10000000_01101011_01110001_10010101_01111011_10000100_01111110_10010011_01100101_01110110_01111111_01101100_01111011_10000101_01110101_01111111_10000101_01111110_10000110_10000000_10001010_10000111_10001101_10000011_01111011_01110001_01100001_10000011_10001010_01110101_10010001_10010110_10000101_01111010_10010101_01111011_01101110_01111011_01101110_10010010_01111001_10000010_01110100_10010000_01110101_10010100_01110011_10001101_10000111_01110001_01111101_10000100_01111001_10000100_01111010_10010010_01111001_10001100;
    //     conv2_bias[95:88] <= 8'b01101011; //normalized bias=107.0000
    //     conv2_weight[13823:12672] <= 1152'b01110111_00110011_10010111_01110110_01000001_10110010_01011010_01110000_10110110_01110110_01110100_10000100_10000010_01101111_10001000_10000010_01111111_10000101_01111011_01111111_01101100_01111001_01111111_10000001_10000100_01101111_10000111_10001111_10000100_10001101_10000011_10000000_10000010_10000011_10000000_01110000_01111010_01101111_10010000_10001001_01111101_01111010_01111111_01111011_10000011_01111110_01101001_01110011_10001010_01110001_01110011_01101000_10010001_01111110_01100110_01111010_10000101_10010111_10000110_10010111_01110101_01110010_01110000_01101011_01110000_01110101_10001100_10001001_10001100_01110100_10001101_10010111_01101110_10000011_10001011_10000111_10000110_01110010_10000010_10010011_10010111_10000101_10000101_10001100_01110001_01111100_10010100_10001011_10000111_10000110_10001001_10000001_10001010_10010110_01110111_10001010_01111000_01100001_10000010_01100011_01111010_01111101_01110111_10001011_10000100_10000111_01111010_01101100_10000101_10000111_10000100_10000001_10001011_10000101_10000011_01011110_10001011_01110100_01110000_10000000_01101001_10010011_01111110_10000000_01110110_01111110_01011011_01111110_10010111_10000101_10001000_01101011_10000000_01111110_10010001_10000100_01101010_01110111_01111100_01101001_10000001_01100101_10011100_10001100;
    //     conv2_bias[103:96] <= 8'b01111100; //normalized bias=124.0000
    //     conv2_weight[14975:13824] <= 1152'b01110000_10010000_01101111_01110101_10000010_01111100_01111010_01110001_01111011_01111101_10000010_10000111_10001011_01110001_01111100_01111110_10000111_01111010_01101001_10001111_01101001_10001000_10000001_10000101_10010100_01101111_01110110_01110100_10001001_10001010_10000011_01111001_10000111_01110111_01110101_10000001_10001101_10000011_01101111_10000000_01111011_10000001_01110000_01110011_01110101_01111100_01101110_01111001_01111011_10001010_01111111_10000110_10100001_10001011_10001010_01110000_01110001_10001000_01100100_01101100_10000001_10000011_10000010_10000010_10000110_10000110_10000000_10001001_10001101_10000111_10010101_01111111_10000101_01101100_10000111_01111101_10010100_10000001_10000101_10011100_01111101_01101010_10001100_01110111_10000000_01110010_01110011_01110000_10011101_10000101_01111111_10001001_01101010_01111010_10000110_10001110_01111011_01110111_10000001_01111101_10001011_10001100_01110100_10010000_10001011_10010000_10010101_01110111_10000100_01110110_01110100_10001100_10010111_01101011_01110000_01111001_01101000_01111000_10001110_10001001_10001110_10010100_01110010_10001100_01111110_10000110_10001111_01110010_01110110_01110001_10001011_10000100_01111011_01110110_01111011_01110000_01110000_01111101_10000000_10011010_10000001_01101000_01111101_10001101;
    //     conv2_bias[111:104] <= 8'b01111110; //normalized bias=126.0000
    //     conv2_weight[16127:14976] <= 1152'b10000010_10010110_10011000_10000000_10100110_10000001_00111100_01001011_01011010_10000111_10000010_01110101_10001010_01111111_10000000_01101100_10001111_01110111_01110011_10001111_01111110_01111111_10000110_01101101_10000000_10000000_01111001_10010000_10000011_10000000_10001010_10000100_01111101_10001000_01111001_01111000_01111010_01111001_10000110_01110000_10000011_10000101_01110101_10001001_01111001_10000101_01110001_10000010_01111010_01111001_10010000_10000101_01110110_01111100_10001111_01110110_01111100_10001011_01111101_01111100_10001100_01111001_10000111_01101111_10001001_10010111_01111100_01111111_01111111_10000011_10000100_10010011_10001001_01111110_01111010_10000100_01101011_10000010_01110110_01111111_01111111_10000010_10001010_01111110_10001001_10000000_10000110_10001100_10000110_01110100_01110100_01101001_01111000_01111011_10000000_01110011_01101011_10010011_10001011_01101101_10000000_01101100_01110010_01100011_10001101_10001000_01110100_10010111_10001010_10000000_10001001_10001001_01111011_10001010_01110010_01101101_01110000_01111001_10001011_01101010_01111010_01110010_10000001_10000001_10001111_10000100_01110110_01110011_01111001_01101010_01110111_10000101_01110100_10000101_01101111_10000110_01111000_10000010_10000110_10001010_10000111_01101111_01110111_01111111;
    //     conv2_bias[119:112] <= 8'b01111111; //normalized bias=127.0000
    //     conv2_weight[17279:16128] <= 1152'b01100110_01110111_01111100_10001100_01100000_01100111_10010000_01101101_01110101_01110110_10001100_01111011_01110101_01110000_10000000_01111111_10000011_01110011_01110011_01111000_10001111_01110010_10000110_10000101_01111011_01101110_01111101_10000111_01111110_10000100_10000011_10000101_01110101_10000111_10001001_01111111_10000000_01111010_10001011_10000101_01111001_10000011_10001001_10010001_01110001_01100110_01111000_10000000_10001110_10001010_01110100_01101110_01110110_10000111_10001001_01110101_01101111_10001010_10001010_01101001_01111110_01111101_10000100_10000100_01110011_10001110_01101110_01111110_01101110_01101001_01111110_01110111_01111111_10000001_10001000_01111101_01110011_10000000_01101101_01110100_01111110_01111101_10001110_10001001_01110010_01111011_10001010_01110110_01110100_10001111_01111101_10000111_01100101_10001011_10000111_01111111_01110001_01111110_10010110_10000101_10000011_10011000_01100010_10001011_10010011_10001101_01111101_01111000_01111010_10000101_10000101_01100100_01100011_10000001_10001010_01110010_10001010_01111101_01110010_01111110_10000111_01111100_10000000_01101110_10000001_10000101_10001000_01111110_10000001_01111101_01111110_10001000_01111011_01110100_01101001_10011001_10000011_10000110_10001010_01110101_10001111_01100101_01111000_10001011;
    //     conv2_bias[127:120] <= 8'b01111011; //normalized bias=123.0000
    //     conv2_weight[18431:17280] <= 1152'b10001111_00111001_10100001_10001110_01010011_10011101_01101110_01011100_10010000_01111010_10010000_01111111_01111000_01110001_01111011_10001111_10001111_10011111_10000100_01110100_01111010_10000111_01111001_01111100_10000010_01111110_10011001_10000100_01110100_10010101_10001101_10010001_01111111_01101010_10001111_01101100_10000110_01111001_01101001_01110001_10000111_10010001_10000000_01110001_01100001_10010000_10000000_01111000_01111101_01110111_10001100_01101111_01111101_01011100_01110101_01110111_10001111_01111001_01011100_01110100_10000101_10001111_01100100_01110111_10000110_01111101_10001101_01110000_10000111_10011010_10001000_10001000_01111000_01111101_10001101_01110100_01111011_10000101_01111101_01111011_01101110_01101000_01111111_01110011_01101001_01110001_01111001_01111001_01110100_01110000_01111110_10001110_10000011_01101111_01110110_10000000_01100111_10010101_10001011_10000101_01101010_10010001_10000011_10001100_01110000_01111000_01110100_01110111_10000110_01111111_01101110_01110000_10010000_01110010_01111010_01110110_10000010_10001000_01111110_01111001_01111111_10000001_10010001_01100101_10001010_10010101_01111110_01100111_01101100_10010001_10001001_01111010_10001111_01110111_01111100_10000011_10001100_01110100_01111101_01110100_10010001_01111110_01110101_01111001;
    //     conv2_bias[135:128] <= 8'b10000100; //normalized bias=132.0000
    //     conv2_weight[19583:18432] <= 1152'b10001001_10100110_10101011_10001011_10001111_10111101_00111111_00100011_01010000_01110011_01111000_10000101_10000011_10001101_10001010_01101110_01111110_01110001_10000001_10000101_01110010_10001101_01111001_01101111_01111101_01111111_10000100_01100111_01101110_01111011_10010101_10000111_10000100_01110110_10001000_01111011_01111111_01101001_01111111_01110010_01111011_10000011_10000000_01111010_01110110_01111011_01111000_10001011_10000000_01111100_10001100_10001000_01110011_10001110_01111111_01111111_01111101_01111010_01111110_10010101_01111000_10000000_01111110_01110101_01011000_10001000_10000101_01101011_01111110_10000010_10000011_01101100_01110001_01110001_01111110_01111110_01111110_01111101_01110111_10000110_10001000_01110000_01110011_01111011_10000010_01101101_10000110_01111100_10000101_10000101_10001110_01110000_10001100_01101110_10001010_01111101_01111111_10000100_10010001_01110100_01100110_10001101_01110110_10010110_01111101_01101101_01110010_10000011_10010000_01101101_01110010_10000100_10001011_01101011_01111011_01100001_10000001_01111110_01110010_10000111_01101100_10000111_01110000_01110010_01110101_10001011_10011000_10000000_10001000_10001010_10000100_01110101_10000101_01111000_10000101_01111000_01111101_10000000_10000010_10000000_01100111_10010011_10000100_01111000;
    //     conv2_bias[143:136] <= 8'b01111100; //normalized bias=124.0000
    //     conv2_weight[20735:19584] <= 1152'b01101000_01101101_01111001_10010101_01100101_01110110_10000111_01001111_10011111_01110110_10000011_01101111_10001010_10000011_01110100_10001010_01110111_01111000_10000000_01111101_10001101_10000001_01101111_10000100_10001011_10001111_10000110_01111110_10000010_01111001_01110100_10000001_10001001_10010000_01110010_10000111_10000010_10010001_01100101_10001001_01101111_10001011_10000001_10001001_10001011_10001000_01111111_01101111_10000100_10100000_10011000_10000100_01111010_01111111_01110010_10000101_10000011_01110010_10010101_10000110_01111111_01111011_10000101_10000001_10010001_10000101_01110110_01110000_01110011_01101011_01110110_10001001_10000101_01101110_10000111_01110111_10000001_01110110_10000100_10001010_10010000_01111101_10000110_10000100_10001000_10000100_01110111_01111011_01110111_01110000_10010010_01111111_10000000_01111111_10001010_01111111_01111111_01111101_01111111_10000100_01101101_10000111_10000100_01110000_10001100_10000010_10000011_10001000_10000111_10001100_10000010_01111100_10010010_10010101_01110010_01100100_10001010_01100010_10000011_01111001_10100000_10010000_10010010_01110011_01110100_01101010_01111100_10001000_01110000_01110010_01101111_01100001_01110000_10001110_01111001_01110111_01101011_10001010_01110101_10001001_01111101_10000000_10001011_01110110;
    //     conv2_bias[151:144] <= 8'b01011101; //normalized bias=93.0000
    //     conv2_weight[21887:20736] <= 1152'b10001111_10001101_01100100_10010100_10100010_00111110_10100110_01111111_01000110_01100011_10010000_10001111_01110110_10011011_10001101_01100011_01111010_10010000_01111101_01101011_01110001_10000110_10010010_01111000_01111001_10000101_01011110_01111001_01111000_10000000_10001101_10001101_10000001_01111010_10001001_10001011_10001001_01111101_01110000_01110001_10001010_10000000_10001110_10001100_01111101_01111110_01111100_01111110_10010010_01111101_01110111_10010110_10000001_01111011_10001010_01101111_10000010_10010001_10001010_01111001_01111010_01110110_01111011_10001111_01111111_01110111_01100110_01111101_01110101_01110011_10001101_10000010_01111100_10001011_10000011_10001001_01110111_01110101_10000000_10001000_01111011_10001100_10001110_10000001_01111001_10001101_01101010_01111010_10001100_01111110_01110011_01110101_01110000_10000111_10000000_01111011_10000010_10000011_10001000_10001010_01110110_01111001_01111101_01111011_10001011_01101101_10011011_01101001_10001000_10001101_10010110_10001110_10000000_01110111_10010001_01111111_01110101_10001101_01101011_10001001_01101110_10000100_01111010_01111010_01111110_10000100_10001000_10000100_10010100_01110100_01110110_10000010_01111110_01110110_01111101_10001011_10000100_01111110_01101000_01110000_10010011_10000000_10011101_10001100;
    //     conv2_bias[159:152] <= 8'b01111101; //normalized bias=125.0000
    //     conv2_weight[23039:21888] <= 1152'b01010111_10001110_01101100_00110110_00001111_01111010_01110110_11001010_10111000_10001001_01111110_01110000_01111011_01110101_01111110_01101101_10000100_01110110_01111010_10010011_01101101_10001010_10000001_10001010_01110111_01111101_01111011_10000010_01100000_01110101_10000111_10000001_01111011_01111111_01111010_10010000_10011100_01110100_01111111_10000011_10000011_01111001_01110011_01110010_01101000_01101001_10001011_10000100_10010011_01111011_10000000_01101110_01101011_01111100_10010011_10000100_10001010_01111000_01110100_10000010_10000000_01110100_01110111_10000111_10000100_01111001_01111101_01101011_01110100_01101001_01111001_01101000_01110000_10000001_10001011_01101101_01111110_01111111_01111011_10001100_10011000_01111010_01110011_01111001_01110010_10010010_10000110_01111101_01110100_01101000_10010100_10000011_10000101_10000100_10000001_01111011_01111110_01111101_01111000_10001101_01111101_01110100_10000110_01110010_01111101_01101110_01111101_10000010_01110111_10001001_10000010_01111010_10001000_01100101_10001000_10001100_01110000_10010000_01101110_01111011_01110110_10000111_01111010_10000010_01110111_01111011_01101111_10000010_01111100_10001011_01110110_01101011_01111111_10000100_10000100_10001101_01111110_01110011_01101000_10001011_01110010_10001000_01101111_10011111;
    //     conv2_bias[167:160] <= 8'b01111100; //normalized bias=124.0000
    //     conv2_weight[24191:23040] <= 1152'b01110111_01000000_10001110_01111001_01100000_10111010_01101010_01011110_10001010_01111101_10000011_10000000_10001111_01101010_10010101_01101010_10001011_10000011_10001000_01101101_10000011_10000010_01101110_10000001_01101111_01110110_10001111_01111001_01110000_10000111_10001001_01101110_10001001_01111010_01110101_01101000_01111010_10000000_01111100_01110010_10001000_10000010_10001000_01110000_10001011_01111000_10001000_01110000_01110111_10001100_01111001_10001110_01101111_01101110_10000001_10000110_01111100_10001110_01111001_10010000_01111011_01110010_01110111_01110001_01101010_01111110_01111111_01111111_10000100_01110000_01111000_01111111_01110101_10000100_10000111_10000000_01110110_10001100_10000010_01111000_10001101_01111100_10000011_01100111_01111101_10001101_01101100_01111000_10010111_01110111_01011101_01110111_01101101_10001011_10010001_10001011_10000011_01110011_01110101_10000111_10000111_10001011_01110001_10001000_01101000_01111011_01111011_01111000_10000010_10010100_01110010_01100111_01111011_10010101_10000010_10010100_10001110_10000101_10000000_01111101_10010011_01110100_01111101_10000101_01101101_01111010_10010000_10001110_01110100_01111111_10010000_01110100_10001010_10000100_10010100_10000111_01111001_01100110_01110110_01111111_10000111_10000010_01111010_01110000;
    //     conv2_bias[175:168] <= 8'b01111010; //normalized bias=122.0000
    //     conv2_weight[25343:24192] <= 1152'b11001100_10011010_10100011_01011000_00110110_01001011_01110011_01110001_10001111_10010011_10000000_10010000_10000110_10000011_10010000_10001001_01111011_10000010_10000011_01111100_01110001_10001011_10001111_10010001_10001110_10001110_10000010_10000001_01100000_10001100_01111011_01101011_10000101_01110000_10001000_10001110_10000001_01101100_01101111_01110000_01110101_10001000_01111110_01110011_10000011_01101111_01111001_01111010_01111100_10001010_10011110_10001110_01101111_01111100_01110010_01111111_10011110_10000100_01111001_10001001_10001010_10000001_10000100_01100111_01111000_10001001_10000010_10010001_01110011_10010010_10011011_01110111_10001011_10001000_01111000_01111000_01100111_10000100_01101111_01110100_01111101_10000001_01111111_10000101_01110111_10000010_01111101_10000011_01111101_10010000_01101100_10000011_10010000_01101111_10000001_01101100_01110100_01111111_01100101_01111011_10001101_10001011_01110100_01110111_01111111_10000111_01111111_01111011_01110101_01111010_10000001_01100111_10000000_01111100_01111001_01111100_01111111_10001111_01111011_01110001_01111011_01110101_01110000_01110010_10000000_10000100_10000001_01100001_01111100_01101101_10010110_01101101_10000011_10000100_01111000_10001011_10000101_01111000_01111110_10001111_01101011_01111011_01111110_10010011;
    //     conv2_bias[183:176] <= 8'b01101011; //normalized bias=107.0000
    //     conv2_weight[26495:25344] <= 1152'b01111110_10011000_01100000_10000100_10010111_01000101_10001000_10101000_01101101_01111100_10010010_10011010_10001011_01101111_01111110_01100011_10000110_10001010_01111000_01110011_10010011_10010111_01111101_10000110_01111110_01101100_01100111_01101100_10000110_10000010_10001100_01110011_01111111_10011100_01111011_01110110_01111000_10001011_01101110_10001101_01111100_01110010_10001010_01101001_01110100_01101110_10010010_10001110_01111110_01111010_01101100_01111111_01110111_01110111_01111100_10001010_01101100_01111100_10000100_01111010_10011100_01111111_01111111_01111000_10011000_10000010_01110000_10011001_01110111_01110010_10011111_01110000_10001011_10100000_10001111_10010100_10000011_10010010_01111000_10001100_10010101_10001001_01110100_10001100_10001001_10000011_10011000_10001010_01101110_01110110_01110011_10001001_10000000_01110101_01101011_10000100_10000000_10000111_01111100_10010011_01111110_01110100_10000100_01111111_10000111_01111101_10100010_10000100_01111100_10010011_10001101_01110001_10001001_01111000_10001010_01110100_10010001_10001100_10001111_01111101_01111100_01110001_01101011_01111001_10000011_10000101_01110100_10001000_01110000_10001000_01101101_10001011_01111000_10001110_01110001_10000001_01111101_01110110_10001100_01111100_10001101_01111100_10001100_01110101;
    //     conv2_bias[191:184] <= 8'b10000110; //normalized bias=134.0000
    //     conv2_weight[27647:26496] <= 1152'b00101010_00001001_00011010_11000100_11100010_10101010_10010110_01111111_10000001_10011001_10000100_01111010_10010011_01111111_10001000_10001000_01111100_10000101_01110010_10000001_10000110_01111111_10000001_01110111_10000100_10010010_10001101_01111100_01110001_01110001_10000001_10001011_01101111_01111101_10000001_01111001_10001000_10011001_10001011_10001010_01111111_10000110_01111110_10100011_10000000_10011011_01110000_10010000_01111101_10001100_10010001_01110100_10000010_10001010_10010001_10000001_10001100_10000001_10010011_01111100_10000110_01111111_10000000_01110101_01111010_10000101_01100111_10000001_01101111_10000001_01110000_10000101_01111010_10000101_01111101_10001010_10000001_01110111_10001101_01111110_10000000_01110111_01111101_01101110_01110111_01110000_10000110_01111010_10001110_01111001_01111111_01110001_10000111_01111001_01110101_10000011_01111101_01111010_10001010_01110011_01110100_01110111_10001010_10001111_01111011_01111101_01111001_01111100_01101111_01110110_10000111_10000010_01101110_10000111_10000011_10010110_01111010_01111011_01111011_01111000_01111100_01101110_01110110_01111100_10010001_10001010_01111010_01111101_01110101_10000001_01111101_01110011_10001001_10010011_10001111_01111000_01111111_01111001_01100010_10000111_10000011_10000000_01110110_10001011;
    //     conv2_bias[199:192] <= 8'b10001000; //normalized bias=136.0000
    //     conv2_weight[28799:27648] <= 1152'b01111001_10100100_10101110_00110011_00011000_01011110_11001111_10001100_10000000_01111101_10001100_10000010_10001110_01111000_10001010_01111101_01111101_01111011_10001101_01111011_10001110_01100000_10000101_10010001_01111001_01111110_01110010_10000110_10010000_10010001_10001001_01111011_01110101_01110000_01100011_01111100_10000011_10001010_01110111_10000111_10010000_01101100_01111101_01110010_10001000_10010011_10000110_01110010_01111110_01110010_10010000_01111101_10000000_10000101_10000101_10000111_01111011_10000010_01110001_10000111_01110010_10000000_01101111_01110011_01111110_01111011_01111100_01101101_01111111_01111100_10000010_10011010_10000010_10001010_10001101_10001110_01101111_10000110_01110010_01100110_01101110_10001100_01111000_01111110_10011000_10010001_01111101_01111010_01111101_01111011_10001100_10000011_01111001_10010101_01110111_01110010_10000010_10000001_10000110_01101101_10000100_01110001_10010011_10000010_10000001_01101100_01111100_01111111_10001010_10001110_10000110_01101100_10000011_10001010_01101100_10001101_01111011_01110001_10000001_01111000_01111001_01111101_01111011_10001000_10000101_10001000_01111100_10000100_01111110_01111000_01111010_10001011_10000010_01111110_10011001_10000001_10000111_10000100_01111101_10000001_10001110_01110110_01111010_01110101;
    //     conv2_bias[207:200] <= 8'b10001010; //normalized bias=138.0000
    //     conv2_weight[29951:28800] <= 1152'b10000111_10000010_10010010_10000001_10100000_10100001_01000101_00111111_01001100_10001010_01110011_01110111_10000010_01110011_01111100_10000101_01111010_10001001_01110101_01110100_10010000_01111110_01110000_01111100_10000001_01111111_10011000_01110101_01110101_01111001_10001101_01101001_01100011_10001110_10001111_01111011_01111001_01100011_10000100_10000001_10000000_01101011_01111100_10001110_01111000_01111111_10000110_01111000_01111011_01111000_01111110_10000110_10000011_01101110_01111011_01111001_10000000_01110111_10010000_01111011_10011100_01111000_01011111_10000110_01111011_10000101_01111010_01111000_01100100_01011100_01111001_10000001_01101111_01110111_01111001_01101001_10000110_10001100_01101011_01111111_10000000_01111011_10000010_01110111_01110001_01110001_01110010_10000100_10010110_01111100_10000010_01111001_10000101_01111110_01111011_10000110_01111100_01110000_01111110_10010101_01110101_01111110_01111000_01111111_01110001_01101111_10000101_10001010_01110000_01110100_01101010_01111111_01110000_01111011_10010000_10000101_10001001_01110010_10010011_10000001_10010010_01111000_01110010_10000010_01101100_10000101_10000100_10010010_10001111_10000111_01110010_01111100_10000000_01110101_01101011_10010011_10000111_01110000_01111001_01111011_10000010_10001110_10000011_01110000;
    //     conv2_bias[215:208] <= 8'b10001110; //normalized bias=142.0000
    //     conv2_weight[31103:29952] <= 1152'b01101001_01100111_01011001_01001111_01101100_01011001_10100011_10011011_10101110_01101110_01101101_10000101_10000001_01101011_10010001_10011001_01100010_10001010_10001010_01101100_10000101_10000001_01110110_10000010_10001010_10001000_01110011_01110000_01111011_01101111_01101101_01110010_10000011_01110011_10000011_10001100_10001110_01110000_10000010_01101010_10001110_01111010_01110001_10001110_10011110_01111011_10001000_10010011_10010111_01110110_01110000_01100000_01111111_01111000_10010101_10000001_01110100_10000011_10010011_10000110_10001000_10011001_10011010_01111011_01101011_01101111_10001010_10000000_10000110_01101110_01011011_10001100_01111010_01110011_01111111_01111111_10000000_01100011_01110010_01100100_01111001_10001010_01111001_10001100_01111111_10001000_01101100_01111101_10000110_01111011_01110111_01111011_01101110_10000111_10001011_01111110_01111001_01111001_01101101_01111010_10000010_01111011_10001000_10000010_10001111_10000001_01111110_01111001_10001001_10001000_01111001_10000101_10001011_01111000_10001100_10000100_01110001_01100111_01111101_10001101_10000101_01100111_10010011_01111101_10001011_10000100_01110010_01110110_10010111_10010001_10000100_01110010_10001001_10010110_01111100_10001100_01111010_01110100_01110110_01111111_10010000_01111000_01101010_10001000;
    //     conv2_bias[223:216] <= 8'b01111110; //normalized bias=126.0000
    //     conv2_weight[32255:31104] <= 1152'b01110101_10000011_01110011_10000000_01111101_01100111_01110111_01110111_01111100_01101110_01100010_10000101_01111110_10000001_01101110_10000101_10010101_10000011_10001100_01111111_10000111_01100111_10000001_10010011_10000011_01110111_01101011_01101011_10000000_01110110_10000001_01111111_10000010_10000011_01100011_10000100_10000110_01110010_01101111_10000011_10001100_01111011_10000100_01111011_01111101_10000100_01110010_01100100_10000011_10000011_01110100_10001100_10001101_10000101_01101000_10000101_01101111_01110000_10010100_10001001_10000010_10001010_10000110_10001010_01110011_01110110_10010010_01110000_01111111_10001100_10000011_10001000_01101101_01111000_01111100_10001001_01110111_01101111_10010111_10000101_10000010_10000010_01111100_01110111_10000010_01111000_10000101_10001000_10001111_01111010_10000000_01111001_01110100_01101010_01111101_01111111_10000001_01111101_01110011_01101100_10010101_01101111_10000000_10000001_10001010_01111011_01101000_10001010_10001110_01101111_01101100_01111111_01110100_10000001_10000101_10001001_10000111_01111010_01111110_01110001_01101101_01111000_10010000_01110001_01111100_01111011_01011111_01110001_01110101_01111001_01110111_01100111_01111010_10001000_01111000_10000100_01110111_10001011_10000010_01111101_01111111_10000011_10010000_01111101;
    //     conv2_bias[231:224] <= 8'b01111101; //normalized bias=125.0000
    //     conv2_weight[33407:32256] <= 1152'b10000110_10001111_10110101_01101111_01000000_01011001_10111010_01101101_01011010_10000010_10011000_01110010_01111001_01111000_10000001_01100011_01101011_01111011_01110101_10000100_10010000_01111000_01111001_01101111_01110100_10000111_10001001_01101000_01110110_10000110_10001110_01111101_01110011_10001000_10000100_10011000_10001101_10000100_01101010_10010010_10011011_10000000_10000110_01101110_10000101_01110000_01110001_10001110_10001100_10000110_10000101_10001010_01110110_10000010_01101100_10000000_01111010_10001110_01110001_10000101_10000001_01110111_01110011_01110111_01100111_10001000_10000011_01111100_10000010_10000000_10000111_10001011_10001000_10000011_01110101_10001010_01101101_01110101_10000000_10010001_01101110_10001011_01111110_10001101_10001001_10000111_10001011_10000000_01111111_01110010_01111110_01111100_01110010_10000110_01111100_10000000_01110111_10000100_01101011_10000100_10010000_01110110_10001100_01101101_01110001_01110000_10001011_01100111_10010111_10000101_01111110_10000000_01110011_10010101_10001001_10000100_10001001_10001010_01111000_10000101_10011011_10010011_01110000_01111100_01110110_10010100_10001110_10010000_01110101_01111100_01110010_01110010_01110000_10000010_01111111_01111010_10001100_01110100_01101111_01100101_01101101_10001100_10001110_10000101;
    //     conv2_bias[239:232] <= 8'b01110100; //normalized bias=116.0000
    //     conv2_weight[34559:33408] <= 1152'b00111001_01001000_01111110_01010001_10111110_10101101_10001001_10101111_01110101_01110111_10000110_01110001_01101010_01110101_10011111_10010110_10000001_01111011_10001000_10000011_10001001_10000101_10000010_01110001_10001110_10000101_01111010_01101010_10000111_01110100_01101100_10001000_10000001_10000010_01101100_01111001_01110000_10001001_01110011_01101011_01110000_01111100_01111111_10000000_10010110_01111011_01111111_10000111_10001110_01101111_10001100_10001001_01110101_01111001_10001000_10010001_01111001_10000000_10011000_01101101_10000111_10011010_10001010_01110111_01110011_01110001_01111101_10001110_10000011_01110111_10001100_01110001_01101100_01110110_01111100_10000001_10000110_10001110_01110000_01100011_01111111_01101111_10000100_10011000_01111110_01101110_01111101_10001000_01110011_10000000_01111100_01111011_10001111_10000110_10001111_10000101_10000010_10001111_01111011_01110100_10010100_10011010_10000101_01110111_01101110_01111111_01111000_10000011_01100100_01101101_10000010_01111000_01111110_10000001_01110101_10000001_01100101_10000001_01111011_10001101_10000010_10001101_01110100_10000010_10010100_10000001_10001111_01111100_10000000_01111100_10000000_01110100_10001101_01110011_01101010_01111010_01101101_10000110_10000011_10001100_01111100_01110011_01110101_01111001;
    //     conv2_bias[247:240] <= 8'b01111000; //normalized bias=120.0000
    //     conv2_weight[35711:34560] <= 1152'b10011100_10111010_10100111_01001011_00101110_00110110_01111000_10100101_10011100_10000010_01111001_10000011_10000100_01110111_01110111_01111100_01111111_10000000_01111111_10001010_10000000_01101001_10000010_10010011_10000011_01110011_10000111_01111001_10001010_01110010_01100111_10000001_01110011_01111001_01110100_01111010_01111010_01110101_01111111_10011100_01111101_10000111_01111110_01101010_10000111_01111100_10000000_01111001_10000100_10010000_10001011_10011101_01110001_10000000_10001110_10001001_01110001_10000110_10000001_01100101_01101101_01111100_01111000_01110010_10001000_10010000_10000010_10010010_01110001_01101110_01110001_10010010_01111101_01101111_01110111_01110010_10000100_10001001_01110111_01101111_10001100_10000110_10000110_10000011_01111101_10001000_01111000_01100111_10011000_10001000_01011001_01111111_01110110_01111111_10000101_10010101_01111000_10001110_01111111_01110001_10000010_01111010_10001101_10000001_01111110_01110100_10000010_10001001_01111000_10011011_01111101_10001100_01111100_10001010_10010011_01111010_10010001_10000010_10000010_01101100_10001011_10000100_10001100_10000110_01101001_01101110_01111111_10000001_01111001_10010000_10000100_01100110_01110001_10000101_01110010_01101111_01101011_01110010_01110010_10001010_10010010_01101110_01110010_10001000;
    //     conv2_bias[255:248] <= 8'b01001010; //normalized bias=74.0000
    //     conv2_weight[36863:35712] <= 1152'b10001001_10010101_10011111_01001011_10001111_10111100_01101101_01101000_10000011_01110100_10001001_01101110_10000010_01110001_10001110_01110111_10010000_01111111_01101101_01101010_10010011_10011110_10000101_10000110_01111100_10100001_01111101_01111111_01101011_10001010_10000000_01111100_01111000_01110110_10001000_01111111_10010010_10000000_10000010_10000011_01111100_10000001_10010110_10010100_01110111_01111011_10000010_10000100_01111110_01110001_10010001_01110100_10000110_10000010_01111010_01111011_01101110_10000000_01100011_01101100_10000010_01111001_01111011_10000010_01101100_01110101_10001001_10000000_01111110_01110000_01110000_10000011_01110000_01111001_10001000_10000110_01110001_10011001_01111010_10001110_01110100_01110100_01110011_01111100_10000010_01101110_10000011_01110101_10000001_01110111_10010000_01111011_10000010_01110000_01111101_10001010_01111110_01110100_10001000_10001110_10000110_10001010_01111001_10010000_01110000_01110110_01111001_01110111_10001111_01111100_10000110_01111111_01110111_01101101_01101101_01111001_01111110_10000100_10010010_01111110_01110101_01110100_01110010_10001001_10001110_10001010_01111101_10001010_01111000_10000110_10000101_10001011_01110111_01101000_10001111_10010111_01110101_10001001_01111111_01111101_10010010_10001100_01111101_01100010;
    // end
endmodule